module Mux2_1(in1, in2, select, data);
	input [31:0] in1, in2, 
	input select;
	output [31:0]data;
	wire [31:0]]andgate1, andgate2, data;
	wire notgate;
	
	genvar i;
	generate
 		for(i=0; i<32; i++) begin : eachMux
 				and a1(andgate1[i], in1[i], select);
				not n1(notgate, select);
				and a2(andgate2[i], in2[i], notgate);
				or o1(data[i], andgate1[i], andgate2[i]);
 	end
 	endgenerate 

endmodule

module Mux2_1_testbench();
	reg in1, in2, select;
	wire data;

	Mux2_1 dut(.in1, .in2, .select, .out);
	initial begin
		select = 0, in1 = 31'b0000 0000 0000 0000 0000 0000 0000 0000 0000 0000 0000 0000 0000 0000 0000 0000, 
		in2 = 31'b0000 0000 0000 0000 0000 0000 0000 0000 0000 0000 0000 0000 0000 0000 0000 0000; #10
		select = 0, in1 = 31'b0000 0000 0000 0000 0000 0000 0000 0000 0000 0000 0000 0000 0000 0000 0000 0000, 
		in2 = 31'b0000 0000 0000 0000 0000 0000 0000 0000 0000 0000 0000 0000 0000 0000 0000 0001; #10
		select = 0, in1 = 31'b0000 0000 0000 0000 0000 0000 0000 0000 0000 0000 0000 0000 0000 0000 0000 0001, 
		in2 = 31'b0000 0000 0000 0000 0000 0000 0000 0000 0000 0000 0000 0000 0000 0000 0000 0000; #10
		select = 0, in1 = 31'b0000 0000 0000 0000 0000 0000 0000 0000 0000 0000 0000 0000 0000 0000 0000 0001, 
		in2 = 31'b0000 0000 0000 0000 0000 0000 0000 0000 0000 0000 0000 0000 0000 0000 0000 0001; #10
		select = 1, in1 = 31'b0000 0000 0000 0000 0000 0000 0000 0000 0000 0000 0000 0000 0000 0000 0000 0000, 
		in2 = 31'b0000 0000 0000 0000 0000 0000 0000 0000 0000 0000 0000 0000 0000 0000 0000 0000; #10
		select = 1, in1 = 31'b0000 0000 0000 0000 0000 0000 0000 0000 0000 0000 0000 0000 0000 0000 0000 0000, 
		in2 = 31'b0000 0000 0000 0000 0000 0000 0000 0000 0000 0000 0000 0000 0000 0000 0000 0001; #10
		select = 1, in1 = 31'b0000 0000 0000 0000 0000 0000 0000 0000 0000 0000 0000 0000 0000 0000 0000 0001, 
		in2 = 31'b0000 0000 0000 0000 0000 0000 0000 0000 0000 0000 0000 0000 0000 0000 0000 0000; #10
		select = 1, in1 = 31'b0000 0000 0000 0000 0000 0000 0000 0000 0000 0000 0000 0000 0000 0000 0000 0001, 
		in2 = 31'b0000 0000 0000 0000 0000 0000 0000 0000 0000 0000 0000 0000 0000 0000 0000 0001; #10
	end
endmodule

